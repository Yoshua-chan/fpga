`timescale 1ns/1ps

module template();

endmodule
